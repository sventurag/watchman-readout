----------------------------------------------------------------------------------
-- Company: IDLAB	
-- Engineer: Salvador Ventura
-- 
-- Create Date: 05/20/2020 10:02:21 PM
-- Design Name:  
-- Module Name: pedestalTrigger - Behavioral
-- Project Name: WATCHMAN
-- Target Devices: MicroZed board
-- Tool Versions: 
-- Description:  Trigger signal to get pedestal arrays
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
 use ieee.numeric_std.all;

entity pedestalTrigger is
    Port ( 
    		clk : in STD_LOGIC;   
           rst : in STD_LOGIC;
           trigger : out STD_LOGIC;   --- output signal 
           mode : in STD_LOGIC;   -- Signal toggling from USER MODE to TRIGGER MODE, 0 for USER MODE, 1 for TRIGGER MODE
           pedestals: in std_logic; -- Signal to start the pedestal acquisition
           average :  in std_logic_vector(31 downto 0); -- Number of averages
           wr_rs:  in std_logic_vector(1 downto 0); -- To synchronize WR and start at window 0
           sstin : in std_logic_vector(2 downto 0)   -- signal for synchronization
           );
end pedestalTrigger;

architecture Behavioral of pedestalTrigger is
type stm_trigger_type is(
   IDLE,
   START,
    WAIT_FOR_NEXT_RUN,
   CNT_START,
   TRIGGER_HIGH_0,
   TRIGGER_LOW_0,
   WAIT_0,
   RUN_NUMBER

   
);

signal stm_trigger : stm_trigger_type := IDLE;
signal cnt_start_i: std_logic_vector(8 downto 0);
signal cnt_intraBuffer_i: std_logic_vector(8 downto 0);
signal cnt_interBuffer_i: std_logic_vector(8 downto 0);
signal cnt_intratrigger : std_logic_vector(13 downto 0);

signal cnt_i : std_logic_vector(8 downto 0);


signal cnt_wait0_i: std_logic_vector(3 downto 0);
signal trigger_i  : std_logic;
signal reg1: std_logic;
signal reg2: std_logic;
signal edge_det_i : std_logic;
signal cnt_average: std_logic_vector(31 downto 0);
signal cnt_run: std_logic_vector(1 downto 0);
signal  wait_number_i: std_logic_vector(3 downto 0);
signal cnt_between_runs_i:  std_logic_vector(26 downto 0);
begin

p_edge_detector :  process(clk)
begin
        if rising_edge (clk) then
            reg1 <= pedestals;
            reg2 <= reg1;
        end if;
   
   
end process p_edge_detector;

edge_det_i <= reg1  and not (reg2);

p_sm:  process(clk,rst, mode ,sstin,pedestals, cnt_run)
  begin 
  
 if (rst = '0') or (mode='0') then
      stm_trigger <= IDLE;
      cnt_start_i <= (others=> '0');
      cnt_i <= (others=> '0');
      cnt_intratrigger<= "10011011111010";
      cnt_wait0_i <= (others=> '0');
            cnt_run <= (others=> '0');
            wait_number_i <=  (others=> '0');
    cnt_between_runs_i<= (others=> '0');
      trigger_i<='0';
      cnt_average<= (others =>'0');
  else 
      if rising_edge(clk) then
          case stm_trigger is
              when IDLE =>
                   if ( edge_det_i= '1')   then 
                       cnt_average<= (others =>'0');                 
                       stm_trigger <= START;
                   else
                       stm_trigger<= IDLE;
                   end if;
               
               when START =>
                            if  (sstin="011")  and (wr_rs="00")  then          -- Sin        
                                      stm_trigger <= CNT_START;
                                       cnt_intratrigger<= "10011011111101";
                              else
                                      stm_trigger<= START;
                                 end if;

              when CNT_START =>
                	   if cnt_start_i <  "000001110" then  -- This synchronization is different for sim and implementation
                   		   	cnt_start_i <= std_logic_vector(unsigned(cnt_start_i) + 1);
           	  	     	   stm_trigger <= CNT_START;           
                 	  else 
                           cnt_start_i <= (others=> '0');
                   		   stm_trigger <= TRIGGER_HIGH_0;
          			 end if;
              when TRIGGER_HIGH_0 =>           
                      trigger_i <= '1';
                      stm_trigger<= TRIGGER_LOW_0;
                      
              when TRIGGER_LOW_0 =>
					   trigger_i <= '0';
	                   if (cnt_intratrigger > "00000000000000" ) then
						  cnt_intratrigger <= std_logic_vector(unsigned(cnt_intratrigger) -1 );
						  stm_trigger <= TRIGGER_LOW_0;
					   else
						  stm_trigger <= RUN_NUMBER;
					   end if;

      when WAIT_0 =>
                        if cnt_wait0_i <= wait_number_i  then
                           cnt_wait0_i <= std_logic_vector(unsigned(cnt_wait0_i) + 1);
                           stm_trigger<= WAIT_0;   
                        else                    
                           stm_trigger <= RUN_NUMBER;
                           cnt_wait0_i<= (others=>'0') ; 
                        end if;
 
     when RUN_NUMBER =>
                        case cnt_run is
                        when "00" =>  -- First RUN over the storage array [ 0,1, 4, 5 ...]
                                    if (cnt_i < "001111111") then    -- First run ends after 128 triggers (one trigger per subBuffer, every subBuffer has 4 windows)
                                       cnt_i <= std_logic_vector(unsigned(cnt_i) + 1);
                                       cnt_intratrigger <= "10011011111101";
                                       stm_trigger <= TRIGGER_HIGH_0;
                                   else
                                         cnt_run <=  std_logic_vector(unsigned(cnt_run) + 1);
                                       stm_trigger <= WAIT_0;
                                       cnt_intratrigger <= "10011011111101";
                                       wait_number_i<="0001";
                                   end if;					  
			           when "01" =>           -- Second RUN over the storage array [1,2, 5, 6...]
                                  if  (cnt_i  < "011111111" ) then   -- Second  run ends after 256 triggers
                                   cnt_i <= std_logic_vector(unsigned(cnt_i) + 1);
                                      cnt_intratrigger <= "10011011111101";
                                      stm_trigger <= TRIGGER_HIGH_0;
                                  else
                                     stm_trigger <= WAIT_0;
                                     cnt_run <=  std_logic_vector(unsigned(cnt_run) + 1);
                                     cnt_intratrigger <= "10011011110101";
                                     wait_number_i<="0001";

                                   end if;
                      
                      when "10" =>           -- Third  RUN over the storage array [2,3,6,7...]
                          if   (cnt_i  < "101111111" ) then  -- Second  run ends after 384  triggers
                               cnt_i <= std_logic_vector(unsigned(cnt_i) + 1);
                               cnt_intratrigger <= "10011011110101";
                               stm_trigger <= TRIGGER_HIGH_0;
                       else
                              stm_trigger <= WAIT_0;
                               cnt_run <=  std_logic_vector(unsigned(cnt_run) + 1);
                               cnt_intratrigger <= "10011011110101";
                                 wait_number_i<="0001";

                        end if;                      
                     
                     when "11" =>     --     Fourth  RUN over the storage array [3,0,7,4,11,8...]
                           if   (cnt_i  <"111111111" ) then  -- Second  run ends after 511  triggers
                                cnt_i <= std_logic_vector(unsigned(cnt_i) + 1);
                                 cnt_intratrigger <= "10011011110101";
                                 stm_trigger <= TRIGGER_HIGH_0;
                             else
                               cnt_i<= (others=>'0') ; 
                                stm_trigger <=WAIT_FOR_NEXT_RUN ;
                                cnt_average<=  std_logic_vector(unsigned(cnt_average) + 1);
                               cnt_run <=  std_logic_vector(unsigned(cnt_run) + 1);
                             end if;
                             
                       when others=> null;
                         end case; 
                         
                          when   WAIT_FOR_NEXT_RUN =>  -- In order to 
                          
                              if cnt_between_runs_i < x"0000010" then -- x"3FFFFF" 
                                    cnt_between_runs_i <= std_logic_vector(unsigned(cnt_between_runs_i) + 1);
                                      stm_trigger<= WAIT_FOR_NEXT_RUN;
                              else
                                       if cnt_average <=average then 
                                         stm_trigger <= START;
                                         cnt_between_runs_i <=(others=>'0');
                                          cnt_start_i <= (others=> '0');

                           else
                                   cnt_start_i <= (others=> '0');
                                   cnt_average<=(others=> '0');
                                   cnt_between_runs_i <=(others=>'0');
                                   stm_trigger<=IDLE;
                                         end if;          
                                end if;

         end case;     
              
     end if;
end if;
          
end process;



trigger<= trigger_i;

end Behavioral;
