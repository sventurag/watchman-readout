---------------------------------------------------------------------------------
-- Company: IDLAB, Hawaii
-- Engineer: Salvador Ventura
-- 
-- Create Date: 09/11/2019
-- Design Name: 
-- Module Name: circularBuffer - 
-- Project Name: WATCHMAN
-- Target Devices: 
-- Tool Versions: 

-- Description: This module controls the writting process in TargetC in function of 
-- a trigger. The main part is done by a state machine with two types of states:
-- hit and wr_add. All the states monitor the trigger signal but the wr_add also
-- contains the logic for moving to the next address. The addresses corresponds to 
-- the number of windows considering 2-windows subbuffers.
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
 use ieee.numeric_std.all;
 use work.TARGETC_pkg.all; --not used in simulations

entity circularBuffer is

 
    port (
    
  clk :            in  std_logic;
  RST :             in  std_logic;  
  trigger :         in std_logic;
  full_fifo :        in std_logic;          
  windowStorage:             in std_logic;
--  enable_write :    out std_logic;
--    enable_write_fifo :    out std_logic;

  RD_add:           out std_logic_vector(8 downto 0);
--  RD_add_fifo:   out std_logic_vector(8 downto 0);
  WR_RS:            out std_logic_vector(1 downto 0);
  WR_CS:            out std_logic_vector(5 downto 0);
  delay_trigger:    in std_logic_vector(3 downto 0);
  Timestamp:        in T_timestamp  -- not used in simulations
  -- Control Signal
 --  CtrlBus_IxSL:    in     T_CtrlBus_IxSL
   
);

end circularBuffer;
 
architecture structure of circularBuffer is
 

COMPONENT rb_output_windowNumber
  PORT (
    clk : IN STD_LOGIC;
    din : IN STD_LOGIC_VECTOR(12 DOWNTO 0);
    wr_en : IN STD_LOGIC;
    rd_en : IN STD_LOGIC;
    dout : OUT STD_LOGIC_VECTOR(12 DOWNTO 0);
    full : OUT STD_LOGIC;
    empty : OUT STD_LOGIC
  );
END COMPONENT;



signal ptr_window_i : std_logic_vector(8 downto 0);
signal counter_i: std_logic_vector(2 downto 0);
signal sstin_i : std_logic;
signal window2read: std_logic_vector(8 downto 0);
signal wr_i: unsigned(8 downto 0);
signal ptr_window_trans_i: std_logic_vector(8 downto 0);
signal fifo_wr_en : std_logic;
signal fifo_rd_en : std_logic;
signal fifo_out: std_logic_vector(12 downto 0);
signal fifo_full : std_logic;
signal fifo_empty: std_logic;
signal flag_number: std_logic_vector(3 downto 0);
signal fifo_out_i: std_logic_vector(12 downto 0);
type stmachine is (start, wr_add ,hit0,hit1, hit2, hit3, hit4, hit5, hit6,hit7,hit8, hit9, hit10, hit11, hit12, hit13,hit14);
signal stm_circularBuffer: stmachine;
signal fifo_in: std_logic_vector(12 downto 0);
signal saved_i: std_logic_vector(8 downto 0);
signal delay_window: std_logic_vector(8 downto 0);
signal  delay_flag : std_logic_vector(3 downto 0);
signal fifo_wr_en_delay: std_logic;
signal current_subBuffer: std_logic_vector(14 downto 0) ;
signal first_round_of_subbuffer: std_logic;
signal jump_wr: std_logic_vector(6 downto 0) ;
signal ptr_window_inter: std_logic_vector(8 downto 0);
signal long_pulse_rst: std_logic;
type stmachine_comp is ( A, B, C, D);

type stmachine_2windows is (retrieve,enable_rd, delay, decide, one_window, two_windowsA, delay2,  two_windowsB);
signal stm_2windows : stmachine_2windows:= enable_rd;
signal enable_write_i: std_logic;
signal cnt_wr_en : std_logic_vector(3 downto 0);
signal cnt_long_pulse : std_logic_vector(3 downto 0);
signal long_pulse_sig: std_logic;
signal trigger_intl: std_logic;
signal rdad_i: std_logic_vector(8 downto 0);
--signal delay_trigger: std_logic_vector(3 downto 0);
attribute mark_debug : string;
type longPulse_type is(
   IDLE,
   LONGPULSE
);

signal longpulse_stm : longpulse_type := IDLE;
attribute mark_debug of window2read: signal is "true";
attribute mark_debug of trigger: signal is "true";
attribute mark_debug of WR_CS: signal is "true";
attribute mark_debug of WR_RS: signal is "true";
attribute mark_debug of wr_i: signal is "true";
attribute mark_debug of ptr_window_i: signal is "true";
attribute fsm_encoding : string;
attribute fsm_encoding of stm_circularBuffer   : signal is "sequential"; 

begin
  ----------------------------------
  -- State machine for handling the trigger and to generate the 
  -- wr/read addresses (signals WR_CS, WR_RS, RD_add and enable_write). 
  
  -- The ptr_window_i counter is running over the number of winwows 
  -- increasing +4 (for a 2-write-address subbuffer).
  
  -- Signal wr_i is ptr_window divided by two (one-bit shift)
  -- to get the real address WR_CS and WR_RS for the TARGETC. This operation
  -- is done in the first state, then, the wr_i is just increased by 1.

  
  -- Signal ptr_sub_i is the current subbuffer window. Uncomment lines were ptr_sub_i appeared
  -- to follow the signal 
  
  -- The first 15 states are for raising flags and to get wr from
  -- the pointer_window_i signal 
  
  
  -- window2read could be modified to get the right window according to the trigger delay
  ----------------------------------
 delay_trigger <= CtrlBus_IxSL.TC_Delay_RB(3 downto 0);

 p_sm:  process(clk,RST, windowStorage,trigger_intl, full_fifo, Timestamp.samplecnt)
variable flag_number_v: std_logic_vector(3 downto 0);
variable current_subBuffer_v: std_logic_vector(14 downto 0) ;
  begin 
 if (RST = '0') or (windowStorage='0') then
      stm_circularBuffer <= start;
      ptr_window_i  <= (others=> '0');
      window2read <= (others=> '0');
      wr_i <= (others=> '0');
      fifo_wr_en <= '0';
      flag_number <= "0000";
      current_subBuffer<= (others=>'0');
      first_round_of_subbuffer <= '1';
      jump_wr<=(others=>'0');

     
  else 
      if rising_edge(clk) then
      case stm_circularBuffer is
      when start =>
           if (windowStorage = '1') and (Timestamp.samplecnt="111") then
           --if (windowStorage = '1') and (counter_i="111") then  -- for simulations only

               stm_circularBuffer <= hit0;
           else
               stm_circularBuffer<= start;
           end if;
         
---------------------------------
-- If a pulse is detected at this point, and taking in account the delay (~8 ns) the pulse ocurred and was sampled in the previous window
---------------------------------    
      when hit0 =>      

          if unsigned(ptr_window_i) /= 0 then
              wr_i <= shift_right(unsigned(ptr_window_i), 1 );  -- Dividing by 2, beacause every WR address in TARGETC corresponds to 2 windows.
            if trigger_intl = '1' then
                flag_number<= "0000";
                window2read <= std_logic_vector(unsigned(ptr_window_i) - 1);
                fifo_wr_en<='1';   
                if  unsigned(delay_trigger)> 0 then 
                 current_subBuffer(0) <='0';
                 jump_wr(0)<= '1';
                else
                 current_subBuffer(0)<='1';
                 jump_wr(0)<= '0';

                end if;   
              
              else
                 fifo_wr_en<='0';  
              end if;
          else
              wr_i <= unsigned(ptr_window_i);
                            
              if trigger_intl = '1' then
                 
                flag_number<= "0000";
                window2read <= std_logic_vector(ptr_window_i);
                fifo_wr_en<='1';   
                 
              else
                 fifo_wr_en<='0';  
              end if;
              
          end if;

          stm_circularBuffer <= hit1;
          
               
          
          

     when hit1 =>      
           if trigger_intl = '1' then
              flag_number<= "0001";

             window2read <= std_logic_vector(ptr_window_i);
             fifo_wr_en<='1';   
             
             if  unsigned(delay_trigger)> 1 then 
                  current_subBuffer(1) <='0';
                  jump_wr(1)<= '1';
             else
                  current_subBuffer(1)<='1';
                  jump_wr(1)<= '0';
             end if;   
           
           else
              fifo_wr_en<='0';    
          end if;
           stm_circularBuffer <= hit2;
 
       
      when hit2 =>      
            if trigger_intl = '1' then
               flag_number<= "0010";

              window2read <= std_logic_vector(ptr_window_i);
              fifo_wr_en<='1';   
              if  unsigned(delay_trigger)> 2 then 
                  current_subBuffer(2) <='0';
                  jump_wr(2)<= '1';
              else
                 current_subBuffer(2)<='1';
                 jump_wr(2)<= '0';
              end if;   
            
              else
               fifo_wr_en<='0';  
           end if;
        stm_circularBuffer <= hit3;
            
---------------------------------
        -- If a pulse is detected at this point, and taking in account the delay (~8 ns) the pulse ocurred and was sampled in the previous window
  ---------------------------------               
       when hit3 =>      
             if trigger_intl = '1' then
                flag_number<= "0011";

              window2read <= std_logic_vector(ptr_window_i);
              fifo_wr_en<='1';   
              if  unsigned(delay_trigger)> 3 then 
                  current_subBuffer(3) <='0';
                  jump_wr(3)<= '1';
              else
                 current_subBuffer(3)<='1';
                 jump_wr(3)<= '0';
              end if;   
             else
--                flag3 <= false;          
                fifo_wr_en<='0';  
                -- window2read <= (others=>'X') ;         
            end if;
           stm_circularBuffer <= hit4;
                     
       
        when hit4 =>      
              if trigger_intl = '1' then
                flag_number<= "0100";

               window2read <= std_logic_vector(unsigned(ptr_window_i) + 1);
               fifo_wr_en<='1';   
              if  unsigned(delay_trigger)> 4 then 
                   current_subBuffer(4) <='0';
                   jump_wr(4)<= '1';
               else
                  current_subBuffer(4)<='1';
                  jump_wr(4)<= '0';
               end if;   
              else
                fifo_wr_en<='0';  
             end if;
           stm_circularBuffer <= hit5;
        
        when hit5 =>      
           if trigger_intl = '1' then
                flag_number<= "0101";

               window2read <= std_logic_vector(unsigned(ptr_window_i) + 1);
               fifo_wr_en<='1';   
              if  unsigned(delay_trigger)> 5 then 
                   current_subBuffer(5) <='0';
                   jump_wr(5)<= '1';
               else
                  current_subBuffer(5)<='1';
                  jump_wr(5)<= '0';
               end if;   
           else
        fifo_wr_en<='0';      
           end if;
             stm_circularBuffer <= hit6;

   
        when hit6 => 
           
           
           ptr_window_inter<= ptr_window_i;
           if trigger_intl = '1' then
                flag_number<= "0110";
              
               window2read <= std_logic_vector(unsigned(ptr_window_i) + 1);
               fifo_wr_en<='1';   
              if  unsigned(delay_trigger)> 6 then 
                   current_subBuffer(6) <='0';
                   jump_wr(6)<= '1';
               else
                  current_subBuffer(6)<='1';
                  jump_wr(6)<= '0';
               end if;   
          else
        fifo_wr_en<='0';  
           end if;
             stm_circularBuffer <= hit7;
             
             
             
       
       when hit7 =>      
        -- In this state, WR and ptr_window are updated,
        --- we have to know if the past states trigger detections
        -- correspond to the first round of the subBuffer, if the 
        -- difference between the delay and the flag is negative (jump_wr)
        -- in order to update WR. 
        -- Suppose the difference is negative, so the trigger  not ocurred in the
        -- current subBuffer, and could correspond to a previous subBuffer
        -- or to the same subBuffer but WR+1
        if first_round_of_subbuffer ='1' then
              if unsigned(ptr_window_i) /=  0 then
                  wr_i <= shift_right(unsigned(ptr_window_i), 1  ) +1;
              else
                  wr_i <= unsigned(ptr_window_i )  + 1 ;
              end if;
                if trigger_intl = '1' then
--                   flag7 <= true;
                    flag_number<= "0111";
                   
                   window2read <= std_logic_vector(unsigned(ptr_window_i) + 1);
                   fifo_wr_en<='1';   
                  if  unsigned(delay_trigger)> 7 then 
                       current_subBuffer(7) <='0';
                   else
                      current_subBuffer(7)<='1';
                   end if;   
               else
                    fifo_wr_en<='0';  
                end if;
                stm_circularBuffer <= hit8;
                jump_wr<=(others=>'0');

              
        else
              if unsigned(jump_wr) > 0 then
                  wr_i <= shift_right(unsigned(ptr_window_i), 1  ) +2;
                  ptr_window_i <=  std_logic_vector(unsigned(ptr_window_inter)+4);
                  jump_wr<=(others=>'0');
                  stm_circularBuffer <= hit0;
 
              else
                  if unsigned(ptr_window_i) /=  0 then
                       wr_i <= shift_right(unsigned(ptr_window_i), 1  ) +1;
                  else
                       wr_i <= unsigned(ptr_window_i )  + 1 ;
                  end if;     
                     if trigger_intl = '1' then
                               flag_number<= "0111";
                              
                              window2read <= std_logic_vector(unsigned(ptr_window_i) + 1);
                              fifo_wr_en<='1';   
                             if  unsigned(delay_trigger)> 7 then 
                                  current_subBuffer(7) <='0';
                              else
                                 current_subBuffer(7)<='1';
                              end if;   
                          else
                               fifo_wr_en<='0';  
                           end if;
                           stm_circularBuffer <= hit8;
                  
               end if;
       end if;           
                                   

  
       when hit8 =>      
             if trigger_intl = '1' then
                flag_number<= "1000";
                
              window2read <= std_logic_vector(unsigned(ptr_window_i) +2); 
              fifo_wr_en<='1';   
              if  unsigned(delay_trigger)> 8 then 
                  current_subBuffer(8) <='0';
              else
                 current_subBuffer(8)<='1';
              end if;       
            else
            fifo_wr_en<='0';  
            end if;
             stm_circularBuffer <= hit9;
           
        when hit9 =>      
              if trigger_intl = '1' then
                flag_number<= "1001";
                 
             window2read <= std_logic_vector(unsigned(ptr_window_i)+2); 
                fifo_wr_en<='1';   
              if  unsigned(delay_trigger)> 9 then 
                    current_subBuffer(9) <='0';
                else
                   current_subBuffer(9)<='1';
                end if;              
              else
                fifo_wr_en<='0';       
             
             end if;
          stm_circularBuffer <= hit10;
          
         when hit10 =>      
               if trigger_intl = '1' then
                flag_number<= "1010";
                  
                  window2read <= std_logic_vector(unsigned(ptr_window_i)+2); 
                fifo_wr_en<='1';   
              if  unsigned(delay_trigger)> 10 then 
                    current_subBuffer(10) <='0';
                else
                   current_subBuffer(10)<='1';
                end if;   
                
               else
              fifo_wr_en<='0';  
              end if;
             stm_circularBuffer <= hit11;
                      
          when hit11 =>      
                if trigger_intl = '1' then
                flag_number<= "1011";
                   
                   window2read <= std_logic_vector(unsigned(ptr_window_i)+2);    
                fifo_wr_en<='1';   
              if  unsigned(delay_trigger)> 11 then 
                    current_subBuffer(11) <='0';
                else
                   current_subBuffer(11)<='1';
                end if;   
                   else
         fifo_wr_en<='0';  
               end if;
             stm_circularBuffer <= hit12;
 
          
          when hit12 =>      
             if trigger_intl = '1' then
                 flag_number<= "1100";
                 window2read <= std_logic_vector(unsigned(ptr_window_i)+3); 
                 fifo_wr_en<='1';   
                 if  unsigned(delay_trigger)> 12 then 
                    current_subBuffer(12) <='0';
                else
                   current_subBuffer(12)<='1';
                end if;   
            else
                   fifo_wr_en<='0';  
            end if;
           
             stm_circularBuffer <= hit13;
  
          when hit13 =>      
             if trigger_intl = '1' then
                flag_number<= "1101";
                 window2read <= std_logic_vector(unsigned(ptr_window_i)+3); 
                fifo_wr_en<='1';   
                
                if  unsigned(delay_trigger)> 13 then 
                    current_subBuffer(13) <='0';
                else
                   current_subBuffer(13)<='1';
                end if;   
             else
                fifo_wr_en<='0';   
             end if;
               stm_circularBuffer <= hit14;             

          when hit14 =>      
             ptr_window_trans_i <= ptr_window_i;
             if trigger_intl = '1' then
             flag_number<= "1110";
                
            window2read <= std_logic_vector(unsigned(ptr_window_i)+3); 
                fifo_wr_en<='1';   
              if  unsigned(delay_trigger)> 14 then 
                    current_subBuffer(14) <='0';
                else
                   current_subBuffer(14)<='1';
                end if;   
             else
                fifo_wr_en<='0';   
      
             end if;
               stm_circularBuffer <= wr_add;
                 
          when wr_add =>
          

          if trigger_intl = '1' then
               flag_number<= "1111";
               window2read <= std_logic_vector(unsigned(ptr_window_i)+3) ; 
               fifo_wr_en<='1';   
               flag_number_v :=flag_number;
               if full_fifo = '0' then
                     if wr_i /= 255 then  
                                ptr_window_i <= std_logic_vector(unsigned(ptr_window_trans_i) + 4);   -- To next subBuffer              
                                 wr_i <= unsigned(wr_i+1);
                                 first_round_of_subbuffer <= '1';
                     else
                          wr_i <= (others => '0');
                     end if;
                     current_subBuffer<= (others=>'0');
     
                   stm_circularBuffer<= hit0;
               else 
                   stm_circularBuffer<= hit0;
               end if;
                             
           else  
                         fifo_wr_en<='0';   
             if  unsigned(current_subBuffer) > 0 then
                 if full_fifo = '0' then

                     ptr_window_i <= std_logic_vector(unsigned(ptr_window_trans_i) + 4);
                     if wr_i /= 255 then  
                         if  unsigned(current_subBuffer) > 0 then           -- To next subBuffer 
                                ptr_window_i <= std_logic_vector(unsigned(ptr_window_trans_i) + 4);                 
        
                               wr_i <= unsigned(wr_i+1); 
                               first_round_of_subbuffer <= '1';
                               long_pulse_rst<='1';
                              else
                               wr_i <= unsigned(wr_i-1);
                               ptr_window_i <= std_logic_vector(unsigned(ptr_window_trans_i) );                 
                               first_round_of_subbuffer <= '0';

                          end if;          
                   
                     else
                               wr_i <= (others => '0');
                     end if;

           
                     stm_circularBuffer<= hit0;
                      current_subBuffer<= (others=>'0');
                 else   
                     stm_circularBuffer<= hit0;  
                      current_subBuffer<= (others=>'0');               
                 end if;
             else  --- NO HIT 
                 current_subBuffer<= (others=>'0');
                 stm_circularBuffer<= hit0;
                 wr_i <= unsigned(wr_i-1);  -- If no hit is detected, the wr pointer goes back to the initial value for the current subBuffer, at this point (the end of wr), 
                                            -- wr - 1 means going back four windows, a subBuffer, so, 
                                            -- the current subBuffer will be overwritted
                first_round_of_subbuffer <= '0';


             end if;             
           stm_circularBuffer <= hit0;
        end if;       
           end case;
   end if;
      
end if;

end process p_sm;
WR_RS <= std_logic_vector(wr_i(1 downto 0));

WR_CS <= std_logic_vector(wr_i(7 downto 2));
----------------------------------
-- Dummy SSTIN signal for simulations
----------------------------------

p_counter: process(clk, RST)
begin
if RST = '0' then
    counter_i <= (others=> '0');
 
else
    if rising_edge(clk) then
        if counter_i < "111" then
           counter_i <= std_logic_vector(unsigned(counter_i) + 1);
        else 
           counter_i <= "000";

        end if;
    end if;
 end if;

end process p_counter;

----------------------------------
-- Dummy signal for simulations
----------------------------------
p_sstin: process(clk,RST)

begin
if RST = '0' then
    sstin_i <= '0';
else
    if rising_edge(clk) then
        case counter_i is 
        when "000" =>
            sstin_i <= '1';
        when "001" =>
            sstin_i <= '1';
        when "010" =>
            sstin_i <= '1';
        when "011" =>
            sstin_i <= '0';
        when "110" => 
           sstin_i <= '0';
        when "111"=> 
           sstin_i <= '1';   
        when others =>
            sstin_i <= '0';
        end case;
     
     end if;
    
 end if;
 

end process p_sstin;

----------------------------------
-- Long pulses handling
----------------------------------
long_pulses_stm:	process(clk,trigger, RST)
       
             
        begin
            if RST = '0' then
                long_pulse_sig <= '0';
                cnt_wr_en <= (others=>'0'); 
      --          trigger_intl<='0';
            else
                if rising_edge(clk) then 
                            case longpulse_stm is
                                 when IDLE =>            
                                if trigger= '1' then           
                                    if cnt_wr_en < "0001" then  --- After x windows (cnt_wr_en < x) the pulse is considered 'long'.
                                        long_pulse_sig<= '0';
                                        cnt_wr_en <= std_logic_vector(unsigned(cnt_wr_en) + 1);
                                        trigger_intl<=trigger;
                                        longpulse_stm <= IDLE;
                                    else
                                        long_pulse_sig<='1';
                                        cnt_wr_en <= (others=>'0');
                                        longpulse_stm <= longpulse;  -- if the writeEn stays high for more than x clk periods the long_pulse signal goes high
                                        trigger_intl<= '0';

                                    end if;    
                               else
                                   long_pulse_sig <= '0';
                                   cnt_wr_en <= (others=>'0');
                                   longpulse_stm <= IDLE;
                                   trigger_intl<=trigger;
                                                
                               end if;
                             when longpulse=>
                                if trigger= '1' then           
                                    long_pulse_sig<= '1';

                                     longpulse_stm <= longpulse; 
                                     trigger_intl<='0';

                                else
                                    long_pulse_sig<= '0';
                                    longpulse_stm <= IDLE;
                                    trigger_intl<=trigger;

                                end if;
                            end case;        
                        
                        end if;
                    end if;
    end process;

----------------------------------
-- Trigger Delay introduced by electronics 
-- For a 4-window subBuffer, a maximum delay of 16 cycles is allowed, as the data is overwritted every 16 cycles
----------------------------------

p_delay_flag : process(clk,RST, delay_trigger,window2read, flag_number)

variable local_window_v:  std_logic_vector(1 downto 0);
variable subtraction_v: integer;
variable delay_flag_v: std_logic_vector(3 downto 0);
variable div_window_v: std_logic_vector(8 downto 0);
begin

if RST = '0' then
    delay_flag_v := (others=> '0');
    delay_window <= (others=> '0');
    local_window_v:=(others=> '0');
    delay_flag <= (others=> '0');
    div_window_v:= (others=> '0');
    
else
    if rising_edge(clk) then 

        div_window_v := std_logic_vector(shift_right(unsigned(window2read), 2  ));
         if unsigned(flag_number) - unsigned(delay_trigger) > 0 then
            delay_flag_v := std_logic_vector(unsigned(flag_number) - unsigned(delay_trigger));
        else
            delay_flag_v := std_logic_vector( 16 + unsigned(flag_number) - unsigned(delay_trigger));
        end if;
        
        case delay_flag_v is
               when "0000" | "0001" | "0010" | "0011" =>
                   local_window_v := "00" ; 
               when "0100" | "0101" | "0110" | "0111" =>
                   local_window_v := "01" ;
               when "1000" | "1001" | "1010" | "1011" =>
                   local_window_v := "10" ;
               when "1100" | "1101" | "1110" | "1111" =>
                   local_window_v := "11" ;
               when others =>
                   local_window_v:= "UU" ;
          end case;
          
         if (unsigned(local_window_v) > unsigned(window2read)) then
            subtraction_v := 4;
         else
            subtraction_v:= 0;
         end if;        
         if unsigned(div_window_v) = 0 then
             delay_window <= "0000000" & local_window_v;
         else
              delay_window <= std_logic_vector(   shift_left(unsigned(div_window_v), 2) - subtraction_v  +   unsigned(local_window_v));    
         end if; 
         delay_flag <=  delay_flag_v;

    end if;
end if;
end process;



p_delay_one_cycle: process(clk,RST, fifo_wr_en)
begin
if RST = '0' then
    fifo_wr_en_delay <= '0';
else
    if rising_edge(clk) then

    fifo_wr_en_delay<= fifo_wr_en;
    end if;
end if;
end process;



fifo_in<= delay_window & delay_flag;


----------------------------------
-- FIFO after RB
----------------------------------
rb_output_windowNumber_inst : rb_output_windowNumber
  PORT MAP (
    clk => clk,
    din => fifo_in,
    wr_en => fifo_wr_en_delay,
    rd_en => fifo_rd_en,
    dout => fifo_out,
    full => fifo_full,
    empty => fifo_empty
  );



----------------------------------
-- One-cycle high for the enable_write 
--- The enable_write is high only once independent of the lenght of the trigger
----------------------------------

p_enableWrite : process(clk,RST)
begin
if RST = '0' then
      saved_i <= (others=> '0');
      enable_write <= '0';

else

    if rising_edge(clk) then
        if rdad_i /= saved_i then
            enable_write <= '1';
            saved_i <= rdad_i;
        else
            enable_write <= '0';
        end if;
     end if;   
end if;

end process p_enableWrite;


----------------------------------
-- one or two windows decision
----------------------------------
p_2window_decision: process(clk,RST)

begin
if RST = '0' then
    rdad_i <= (others=> '0');
    enable_write_i <= '0';
    fifo_rd_en <= '0';
    fifo_out_i <= (others=> '0');
else    
    if rising_edge(clk) then 
        case stm_2windows is
            when enable_rd =>
                enable_write_i <= '0';
                if fifo_empty = '0' then
                      fifo_rd_en <= '1';
                      stm_2windows <=delay;
                else 
                    stm_2windows <= enable_rd;
                end if;
             
            when delay=>
                 fifo_rd_en <= '0';
                enable_write_i <= '0';
                  stm_2windows <=retrieve ;
           when retrieve =>
            fifo_out_i <= fifo_out;
            stm_2windows <=decide;
          
            when decide =>
                  fifo_rd_en <= '0';                
                case fifo_out_i(3 downto 0) is -- flag numbers
                    when "0011" | "0111" |"1011" => -- FIX '0000' case not handled 
                    stm_2windows <= two_windowsA;
                    when others =>
                    stm_2windows <= one_window;
                end case;
                enable_write_i <= '0';
                
            when two_windowsA=>
                rdad_i <=   fifo_out_i(12 downto 4);
                enable_write_i <= '1';
                stm_2windows <= delay2;
          
            when delay2=>
                     fifo_rd_en <= '0';
                    enable_write_i <= '0';
                      stm_2windows <=two_windowsB ;
                      
            when two_windowsB=>
                    rdad_i <=std_logic_vector(unsigned(fifo_out_i(12 downto 4)) +1); 
                    enable_write_i <= '1';
                    stm_2windows <= enable_rd;
                    

            when one_window=>
                rdad_i <= fifo_out_i(12 downto 4);
                enable_write_i <= '1';
                stm_2windows <= enable_rd;
    
           end case;
    end if;
end if;
end process;




end architecture;